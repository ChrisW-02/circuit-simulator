* A purely resistive circuit with AC current sources
R1 N001 0 4
R2 N002 0 6
R3 N003 0 8
R4 N002 N001 3
R5 N003 N002 5
R6 N003 N001 6
I1 0 N001 AC(6 0)
I2 N001 N003 AC(4 0)
.ac dec 10 100 10k 
.end