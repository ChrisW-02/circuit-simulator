I1 0 N001 AC(3 0)
R1 N001 N002 5
R2 0 N002 10
R3 N002 N003 20
R4 0 N003 5
R5 0 N004 2
I2 N003 N004 AC(7 0)
.ac dec 10 10 100k
.end
